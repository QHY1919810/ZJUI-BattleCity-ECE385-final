module randomgenerate(input logic Clk ,output logic [30:0]o);   //(2*5)*4
    xor (t0,o[0],o[1]);
    assign t1=o[0];
    assign t2=o[1];
    assign t3=o[2];
    assign t4=o[3];
	 assign t5=o[4];
    assign t6=o[5];
    assign t7=o[6];
    assign t8=o[7];
	 assign t9=o[8];
	 assign t10=o[9];
    assign t11=o[10];
    assign t12=o[11];
    assign t13=o[12];
	 assign t14=o[13];
    assign t15=o[14];
    assign t16=o[15];
    assign t17=o[16];
	 assign t18=o[17];
	 assign t19=o[18];
	 assign t20=o[19];
    assign t21=o[20];
    assign t22=o[21];
    assign t23=o[22];
	 assign t24=o[23];
    assign t25=o[24];
    assign t26=o[25];
    assign t27=o[26];
	 assign t28=o[27];
	 assign t29=o[28];
	 assign t30=o[29];
    assign t31=o[30];
    tff0 u1(.q(o[0]),.t(t0),.c(Clk));
    tff1 u2(.q(o[1]),.t(t1),.c(Clk));
    tff1 u3(.q(o[2]),.t(t2),.c(Clk));
    tff1 u4(.q(o[3]),.t(t3),.c(Clk));
    tff1 u5(.q(o[4]),.t(t4),.c(Clk));
	 tff1 u6(.q(o[5]),.t(t5),.c(Clk));
	 tff1 u7(.q(o[6]),.t(t6),.c(Clk));
	 tff1 u8(.q(o[7]),.t(t7),.c(Clk));
	 tff1 u9(.q(o[8]),.t(t8),.c(Clk));
	 tff1 u10(.q(o[9]),.t(t9),.c(Clk));
	 tff1 u11(.q(o[10]),.t(t10),.c(Clk));
    tff1 u12(.q(o[11]),.t(t11),.c(Clk));
    tff1 u13(.q(o[12]),.t(t12),.c(Clk));
    tff1 u14(.q(o[13]),.t(t13),.c(Clk));
    tff1 u15(.q(o[14]),.t(t14),.c(Clk));
	 tff1 u16(.q(o[15]),.t(t15),.c(Clk));
	 tff1 u17(.q(o[16]),.t(t16),.c(Clk));
	 tff1 u18(.q(o[17]),.t(t17),.c(Clk));
	 tff1 u19(.q(o[18]),.t(t18),.c(Clk));
	 tff1 u20(.q(o[19]),.t(t19),.c(Clk));
	 tff1 u21(.q(o[20]),.t(t20),.c(Clk));
    tff1 u22(.q(o[21]),.t(t21),.c(Clk));
    tff1 u23(.q(o[22]),.t(t22),.c(Clk));
    tff1 u24(.q(o[23]),.t(t23),.c(Clk));
    tff1 u25(.q(o[24]),.t(t24),.c(Clk));
	 tff1 u26(.q(o[25]),.t(t25),.c(Clk));
	 tff1 u27(.q(o[26]),.t(t26),.c(Clk));
	 tff1 u28(.q(o[27]),.t(t27),.c(Clk));
	 tff1 u29(.q(o[28]),.t(t28),.c(Clk));
	 tff1 u30(.q(o[29]),.t(t29),.c(Clk));
	 tff1 u31(.q(o[30]),.t(t30),.c(Clk));
	 
endmodule